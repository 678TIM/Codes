// Code your design here
`include "top.sv"
`include "mips.sv"
`include "imem.sv"
`include "dmem.sv"
`include "controller.sv"
`include "datapath.sv"
`include "maindec.sv"
`include "aludec.sv"
`include "flopr.sv"
`include "adder.sv"
`include "sl2.sv"
`include "mux2.sv"
`include "0706_regfile.sv"
`include "signext.sv"
`include "alu.sv"
`include "sl16.sv"
`include "mux4.sv"
`include "zeroext.sv"